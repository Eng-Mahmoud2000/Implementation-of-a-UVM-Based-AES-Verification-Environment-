package pack1;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "sequence_item_class.sv"
    `include "sequence_class.sv"
    `include "sequencer_class.sv"
    `include "driver_class.sv"
    `include "monitor_class.sv"
    `include "subscriber_class.sv"
    `include "scoreboard_class.sv"
    `include "agent_class.sv"
    `include "env_class.sv"
    `include "test_class.sv"
endpackage




  