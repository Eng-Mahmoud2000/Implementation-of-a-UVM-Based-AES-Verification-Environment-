interface intf();
// input & output signals
logic       [127:0] Data_in;
logic       [127:0] key;
logic       [127:0] Data_out;

endinterface

  